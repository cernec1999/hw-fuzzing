module lock(
    input wire reset_n,
    input wire clk,

    input wire [3:0] code,
    output wire [5:0] state,
    output wire unlocked
    );

    reg [5:0] __reg_state_0;
    wire [5:0] __reg_state_0_next;

    always @(posedge clk, negedge reset_n) begin
        if (~reset_n) begin
            __reg_state_0 <= 6'h0;
        end
        else begin
            __reg_state_0 <= __reg_state_0_next;
        end
    end

    wire __temp_0;
    wire __temp_1;
    wire __temp_2;
    wire __temp_3;
    wire [5:0] __temp_4;
    wire __temp_5;
    wire __temp_6;
    wire __temp_7;
    wire [5:0] __temp_8;
    wire __temp_9;
    wire __temp_10;
    wire __temp_11;
    wire [5:0] __temp_12;
    wire __temp_13;
    wire __temp_14;
    wire __temp_15;
    wire [5:0] __temp_16;
    wire __temp_17;
    wire __temp_18;
    wire __temp_19;
    wire [5:0] __temp_20;
    wire __temp_21;
    wire __temp_22;
    wire __temp_23;
    wire [5:0] __temp_24;
    wire __temp_25;
    wire __temp_26;
    wire __temp_27;
    wire [5:0] __temp_28;
    wire __temp_29;
    wire __temp_30;
    wire __temp_31;
    wire [5:0] __temp_32;
    wire __temp_33;
    wire __temp_34;
    wire __temp_35;
    wire [5:0] __temp_36;
    wire __temp_37;
    wire __temp_38;
    wire __temp_39;
    wire [5:0] __temp_40;
    wire __temp_41;
    wire __temp_42;
    wire __temp_43;
    wire [5:0] __temp_44;
    wire __temp_45;
    wire __temp_46;
    wire __temp_47;
    wire [5:0] __temp_48;
    wire __temp_49;
    wire __temp_50;
    wire __temp_51;
    wire [5:0] __temp_52;
    wire __temp_53;
    wire __temp_54;
    wire __temp_55;
    wire [5:0] __temp_56;
    wire __temp_57;
    wire __temp_58;
    wire __temp_59;
    wire [5:0] __temp_60;
    wire __temp_61;
    wire __temp_62;
    wire __temp_63;
    wire [5:0] __temp_64;
    wire __temp_65;
    wire __temp_66;
    wire __temp_67;
    wire [5:0] __temp_68;
    wire __temp_69;
    wire __temp_70;
    wire __temp_71;
    wire [5:0] __temp_72;
    wire __temp_73;
    wire __temp_74;
    wire __temp_75;
    wire [5:0] __temp_76;
    wire __temp_77;
    wire __temp_78;
    wire __temp_79;
    wire [5:0] __temp_80;
    wire __temp_81;
    wire __temp_82;
    wire __temp_83;
    wire [5:0] __temp_84;
    wire __temp_85;
    wire __temp_86;
    wire __temp_87;
    wire [5:0] __temp_88;
    wire __temp_89;
    wire __temp_90;
    wire __temp_91;
    wire [5:0] __temp_92;
    wire __temp_93;
    wire __temp_94;
    wire __temp_95;
    wire [5:0] __temp_96;
    wire __temp_97;
    wire __temp_98;
    wire __temp_99;
    wire [5:0] __temp_100;
    wire __temp_101;
    wire __temp_102;
    wire __temp_103;
    wire [5:0] __temp_104;
    wire __temp_105;
    wire __temp_106;
    wire __temp_107;
    wire [5:0] __temp_108;
    wire __temp_109;
    wire __temp_110;
    wire __temp_111;
    wire [5:0] __temp_112;
    wire __temp_113;
    wire __temp_114;
    wire __temp_115;
    wire [5:0] __temp_116;
    wire __temp_117;
    wire __temp_118;
    wire __temp_119;
    wire [5:0] __temp_120;
    wire __temp_121;
    wire __temp_122;
    wire __temp_123;
    wire [5:0] __temp_124;
    wire __temp_125;
    wire __temp_126;
    wire __temp_127;
    wire [5:0] __temp_128;
    wire __temp_129;
    wire __temp_130;
    wire __temp_131;
    wire [5:0] __temp_132;
    wire __temp_133;
    wire __temp_134;
    wire __temp_135;
    wire [5:0] __temp_136;
    wire __temp_137;
    wire __temp_138;
    wire __temp_139;
    wire [5:0] __temp_140;
    wire __temp_141;
    wire __temp_142;
    wire __temp_143;
    wire [5:0] __temp_144;
    wire __temp_145;
    wire __temp_146;
    wire __temp_147;
    wire [5:0] __temp_148;
    wire __temp_149;
    wire __temp_150;
    wire __temp_151;
    wire [5:0] __temp_152;
    wire __temp_153;
    wire __temp_154;
    wire __temp_155;
    wire [5:0] __temp_156;
    wire __temp_157;
    wire __temp_158;
    wire __temp_159;
    wire [5:0] __temp_160;
    wire __temp_161;
    wire __temp_162;
    wire __temp_163;
    wire [5:0] __temp_164;
    wire __temp_165;
    wire __temp_166;
    wire __temp_167;
    wire [5:0] __temp_168;
    wire __temp_169;
    wire __temp_170;
    wire __temp_171;
    wire [5:0] __temp_172;
    wire __temp_173;
    wire __temp_174;
    wire __temp_175;
    wire [5:0] __temp_176;
    wire __temp_177;
    wire __temp_178;
    wire __temp_179;
    wire [5:0] __temp_180;
    wire __temp_181;
    wire __temp_182;
    wire __temp_183;
    wire [5:0] __temp_184;
    wire __temp_185;
    wire __temp_186;
    wire __temp_187;
    wire [5:0] __temp_188;
    wire __temp_189;
    wire __temp_190;
    wire __temp_191;
    wire [5:0] __temp_192;
    wire __temp_193;
    wire __temp_194;
    wire __temp_195;
    wire [5:0] __temp_196;
    wire __temp_197;
    wire __temp_198;
    wire __temp_199;
    wire [5:0] __temp_200;
    wire __temp_201;
    wire __temp_202;
    wire __temp_203;
    wire [5:0] __temp_204;
    wire __temp_205;
    wire __temp_206;
    wire __temp_207;
    wire [5:0] __temp_208;
    wire __temp_209;
    wire __temp_210;
    wire __temp_211;
    wire [5:0] __temp_212;
    wire __temp_213;
    wire __temp_214;
    wire __temp_215;
    wire [5:0] __temp_216;
    wire __temp_217;
    wire __temp_218;
    wire __temp_219;
    wire [5:0] __temp_220;
    wire __temp_221;
    wire __temp_222;
    wire __temp_223;
    wire [5:0] __temp_224;
    wire __temp_225;
    wire __temp_226;
    wire __temp_227;
    wire [5:0] __temp_228;
    wire __temp_229;
    wire __temp_230;
    wire __temp_231;
    wire [5:0] __temp_232;
    wire __temp_233;
    wire __temp_234;
    wire __temp_235;
    wire [5:0] __temp_236;
    wire __temp_237;
    wire __temp_238;
    wire __temp_239;
    wire [5:0] __temp_240;
    wire __temp_241;
    wire __temp_242;
    wire __temp_243;
    wire [5:0] __temp_244;
    wire __temp_245;
    wire __temp_246;
    wire __temp_247;
    wire [5:0] __temp_248;
    wire __temp_249;
    wire __temp_250;
    wire __temp_251;
    wire [5:0] __temp_252;

    assign state = __reg_state_0;
    assign __temp_0 = __reg_state_0 == 6'h3f;
    assign unlocked = __temp_0;
    assign __temp_1 = code == 4'h8;
    assign __temp_2 = __reg_state_0 == 6'h0;
    assign __temp_3 = __temp_2 & __temp_1;
    assign __temp_4 = __temp_3 ? 6'h1 : __reg_state_0;
    assign __temp_5 = code == 4'hf;
    assign __temp_6 = __reg_state_0 == 6'h1;
    assign __temp_7 = __temp_6 & __temp_5;
    assign __temp_8 = __temp_7 ? 6'h2 : __temp_4;
    assign __temp_9 = code == 4'h2;
    assign __temp_10 = __reg_state_0 == 6'h2;
    assign __temp_11 = __temp_10 & __temp_9;
    assign __temp_12 = __temp_11 ? 6'h3 : __temp_8;
    assign __temp_13 = code == 4'h7;
    assign __temp_14 = __reg_state_0 == 6'h3;
    assign __temp_15 = __temp_14 & __temp_13;
    assign __temp_16 = __temp_15 ? 6'h4 : __temp_12;
    assign __temp_17 = code == 4'h1;
    assign __temp_18 = __reg_state_0 == 6'h4;
    assign __temp_19 = __temp_18 & __temp_17;
    assign __temp_20 = __temp_19 ? 6'h5 : __temp_16;
    assign __temp_21 = code == 4'hd;
    assign __temp_22 = __reg_state_0 == 6'h5;
    assign __temp_23 = __temp_22 & __temp_21;
    assign __temp_24 = __temp_23 ? 6'h6 : __temp_20;
    assign __temp_25 = code == 4'he;
    assign __temp_26 = __reg_state_0 == 6'h6;
    assign __temp_27 = __temp_26 & __temp_25;
    assign __temp_28 = __temp_27 ? 6'h7 : __temp_24;
    assign __temp_29 = code == 4'h7;
    assign __temp_30 = __reg_state_0 == 6'h7;
    assign __temp_31 = __temp_30 & __temp_29;
    assign __temp_32 = __temp_31 ? 6'h8 : __temp_28;
    assign __temp_33 = code == 4'h9;
    assign __temp_34 = __reg_state_0 == 6'h8;
    assign __temp_35 = __temp_34 & __temp_33;
    assign __temp_36 = __temp_35 ? 6'h9 : __temp_32;
    assign __temp_37 = code == 4'h8;
    assign __temp_38 = __reg_state_0 == 6'h9;
    assign __temp_39 = __temp_38 & __temp_37;
    assign __temp_40 = __temp_39 ? 6'ha : __temp_36;
    assign __temp_41 = code == 4'hb;
    assign __temp_42 = __reg_state_0 == 6'ha;
    assign __temp_43 = __temp_42 & __temp_41;
    assign __temp_44 = __temp_43 ? 6'hb : __temp_40;
    assign __temp_45 = code == 4'h6;
    assign __temp_46 = __reg_state_0 == 6'hb;
    assign __temp_47 = __temp_46 & __temp_45;
    assign __temp_48 = __temp_47 ? 6'hc : __temp_44;
    assign __temp_49 = code == 4'he;
    assign __temp_50 = __reg_state_0 == 6'hc;
    assign __temp_51 = __temp_50 & __temp_49;
    assign __temp_52 = __temp_51 ? 6'hd : __temp_48;
    assign __temp_53 = code == 4'he;
    assign __temp_54 = __reg_state_0 == 6'hd;
    assign __temp_55 = __temp_54 & __temp_53;
    assign __temp_56 = __temp_55 ? 6'he : __temp_52;
    assign __temp_57 = code == 4'h1;
    assign __temp_58 = __reg_state_0 == 6'he;
    assign __temp_59 = __temp_58 & __temp_57;
    assign __temp_60 = __temp_59 ? 6'hf : __temp_56;
    assign __temp_61 = code == 4'h1;
    assign __temp_62 = __reg_state_0 == 6'hf;
    assign __temp_63 = __temp_62 & __temp_61;
    assign __temp_64 = __temp_63 ? 6'h10 : __temp_60;
    assign __temp_65 = code == 4'h5;
    assign __temp_66 = __reg_state_0 == 6'h10;
    assign __temp_67 = __temp_66 & __temp_65;
    assign __temp_68 = __temp_67 ? 6'h11 : __temp_64;
    assign __temp_69 = code == 4'he;
    assign __temp_70 = __reg_state_0 == 6'h11;
    assign __temp_71 = __temp_70 & __temp_69;
    assign __temp_72 = __temp_71 ? 6'h12 : __temp_68;
    assign __temp_73 = code == 4'h9;
    assign __temp_74 = __reg_state_0 == 6'h12;
    assign __temp_75 = __temp_74 & __temp_73;
    assign __temp_76 = __temp_75 ? 6'h13 : __temp_72;
    assign __temp_77 = code == 4'h7;
    assign __temp_78 = __reg_state_0 == 6'h13;
    assign __temp_79 = __temp_78 & __temp_77;
    assign __temp_80 = __temp_79 ? 6'h14 : __temp_76;
    assign __temp_81 = code == 4'hf;
    assign __temp_82 = __reg_state_0 == 6'h14;
    assign __temp_83 = __temp_82 & __temp_81;
    assign __temp_84 = __temp_83 ? 6'h15 : __temp_80;
    assign __temp_85 = code == 4'hf;
    assign __temp_86 = __reg_state_0 == 6'h15;
    assign __temp_87 = __temp_86 & __temp_85;
    assign __temp_88 = __temp_87 ? 6'h16 : __temp_84;
    assign __temp_89 = code == 4'h4;
    assign __temp_90 = __reg_state_0 == 6'h16;
    assign __temp_91 = __temp_90 & __temp_89;
    assign __temp_92 = __temp_91 ? 6'h17 : __temp_88;
    assign __temp_93 = code == 4'h5;
    assign __temp_94 = __reg_state_0 == 6'h17;
    assign __temp_95 = __temp_94 & __temp_93;
    assign __temp_96 = __temp_95 ? 6'h18 : __temp_92;
    assign __temp_97 = code == 4'hf;
    assign __temp_98 = __reg_state_0 == 6'h18;
    assign __temp_99 = __temp_98 & __temp_97;
    assign __temp_100 = __temp_99 ? 6'h19 : __temp_96;
    assign __temp_101 = code == 4'hc;
    assign __temp_102 = __reg_state_0 == 6'h19;
    assign __temp_103 = __temp_102 & __temp_101;
    assign __temp_104 = __temp_103 ? 6'h1a : __temp_100;
    assign __temp_105 = code == 4'h1;
    assign __temp_106 = __reg_state_0 == 6'h1a;
    assign __temp_107 = __temp_106 & __temp_105;
    assign __temp_108 = __temp_107 ? 6'h1b : __temp_104;
    assign __temp_109 = code == 4'ha;
    assign __temp_110 = __reg_state_0 == 6'h1b;
    assign __temp_111 = __temp_110 & __temp_109;
    assign __temp_112 = __temp_111 ? 6'h1c : __temp_108;
    assign __temp_113 = code == 4'h1;
    assign __temp_114 = __reg_state_0 == 6'h1c;
    assign __temp_115 = __temp_114 & __temp_113;
    assign __temp_116 = __temp_115 ? 6'h1d : __temp_112;
    assign __temp_117 = code == 4'h8;
    assign __temp_118 = __reg_state_0 == 6'h1d;
    assign __temp_119 = __temp_118 & __temp_117;
    assign __temp_120 = __temp_119 ? 6'h1e : __temp_116;
    assign __temp_121 = code == 4'h8;
    assign __temp_122 = __reg_state_0 == 6'h1e;
    assign __temp_123 = __temp_122 & __temp_121;
    assign __temp_124 = __temp_123 ? 6'h1f : __temp_120;
    assign __temp_125 = code == 4'h5;
    assign __temp_126 = __reg_state_0 == 6'h1f;
    assign __temp_127 = __temp_126 & __temp_125;
    assign __temp_128 = __temp_127 ? 6'h20 : __temp_124;
    assign __temp_129 = code == 4'h4;
    assign __temp_130 = __reg_state_0 == 6'h20;
    assign __temp_131 = __temp_130 & __temp_129;
    assign __temp_132 = __temp_131 ? 6'h21 : __temp_128;
    assign __temp_133 = code == 4'h9;
    assign __temp_134 = __reg_state_0 == 6'h21;
    assign __temp_135 = __temp_134 & __temp_133;
    assign __temp_136 = __temp_135 ? 6'h22 : __temp_132;
    assign __temp_137 = code == 4'he;
    assign __temp_138 = __reg_state_0 == 6'h22;
    assign __temp_139 = __temp_138 & __temp_137;
    assign __temp_140 = __temp_139 ? 6'h23 : __temp_136;
    assign __temp_141 = code == 4'hc;
    assign __temp_142 = __reg_state_0 == 6'h23;
    assign __temp_143 = __temp_142 & __temp_141;
    assign __temp_144 = __temp_143 ? 6'h24 : __temp_140;
    assign __temp_145 = code == 4'h1;
    assign __temp_146 = __reg_state_0 == 6'h24;
    assign __temp_147 = __temp_146 & __temp_145;
    assign __temp_148 = __temp_147 ? 6'h25 : __temp_144;
    assign __temp_149 = code == 4'h9;
    assign __temp_150 = __reg_state_0 == 6'h25;
    assign __temp_151 = __temp_150 & __temp_149;
    assign __temp_152 = __temp_151 ? 6'h26 : __temp_148;
    assign __temp_153 = code == 4'hf;
    assign __temp_154 = __reg_state_0 == 6'h26;
    assign __temp_155 = __temp_154 & __temp_153;
    assign __temp_156 = __temp_155 ? 6'h27 : __temp_152;
    assign __temp_157 = code == 4'h5;
    assign __temp_158 = __reg_state_0 == 6'h27;
    assign __temp_159 = __temp_158 & __temp_157;
    assign __temp_160 = __temp_159 ? 6'h28 : __temp_156;
    assign __temp_161 = code == 4'h6;
    assign __temp_162 = __reg_state_0 == 6'h28;
    assign __temp_163 = __temp_162 & __temp_161;
    assign __temp_164 = __temp_163 ? 6'h29 : __temp_160;
    assign __temp_165 = code == 4'he;
    assign __temp_166 = __reg_state_0 == 6'h29;
    assign __temp_167 = __temp_166 & __temp_165;
    assign __temp_168 = __temp_167 ? 6'h2a : __temp_164;
    assign __temp_169 = code == 4'h5;
    assign __temp_170 = __reg_state_0 == 6'h2a;
    assign __temp_171 = __temp_170 & __temp_169;
    assign __temp_172 = __temp_171 ? 6'h2b : __temp_168;
    assign __temp_173 = code == 4'h9;
    assign __temp_174 = __reg_state_0 == 6'h2b;
    assign __temp_175 = __temp_174 & __temp_173;
    assign __temp_176 = __temp_175 ? 6'h2c : __temp_172;
    assign __temp_177 = code == 4'h4;
    assign __temp_178 = __reg_state_0 == 6'h2c;
    assign __temp_179 = __temp_178 & __temp_177;
    assign __temp_180 = __temp_179 ? 6'h2d : __temp_176;
    assign __temp_181 = code == 4'h8;
    assign __temp_182 = __reg_state_0 == 6'h2d;
    assign __temp_183 = __temp_182 & __temp_181;
    assign __temp_184 = __temp_183 ? 6'h2e : __temp_180;
    assign __temp_185 = code == 4'h9;
    assign __temp_186 = __reg_state_0 == 6'h2e;
    assign __temp_187 = __temp_186 & __temp_185;
    assign __temp_188 = __temp_187 ? 6'h2f : __temp_184;
    assign __temp_189 = code == 4'hc;
    assign __temp_190 = __reg_state_0 == 6'h2f;
    assign __temp_191 = __temp_190 & __temp_189;
    assign __temp_192 = __temp_191 ? 6'h30 : __temp_188;
    assign __temp_193 = code == 4'hb;
    assign __temp_194 = __reg_state_0 == 6'h30;
    assign __temp_195 = __temp_194 & __temp_193;
    assign __temp_196 = __temp_195 ? 6'h31 : __temp_192;
    assign __temp_197 = code == 4'h6;
    assign __temp_198 = __reg_state_0 == 6'h31;
    assign __temp_199 = __temp_198 & __temp_197;
    assign __temp_200 = __temp_199 ? 6'h32 : __temp_196;
    assign __temp_201 = code == 4'h4;
    assign __temp_202 = __reg_state_0 == 6'h32;
    assign __temp_203 = __temp_202 & __temp_201;
    assign __temp_204 = __temp_203 ? 6'h33 : __temp_200;
    assign __temp_205 = code == 4'h3;
    assign __temp_206 = __reg_state_0 == 6'h33;
    assign __temp_207 = __temp_206 & __temp_205;
    assign __temp_208 = __temp_207 ? 6'h34 : __temp_204;
    assign __temp_209 = code == 4'h8;
    assign __temp_210 = __reg_state_0 == 6'h34;
    assign __temp_211 = __temp_210 & __temp_209;
    assign __temp_212 = __temp_211 ? 6'h35 : __temp_208;
    assign __temp_213 = code == 4'h4;
    assign __temp_214 = __reg_state_0 == 6'h35;
    assign __temp_215 = __temp_214 & __temp_213;
    assign __temp_216 = __temp_215 ? 6'h36 : __temp_212;
    assign __temp_217 = code == 4'hc;
    assign __temp_218 = __reg_state_0 == 6'h36;
    assign __temp_219 = __temp_218 & __temp_217;
    assign __temp_220 = __temp_219 ? 6'h37 : __temp_216;
    assign __temp_221 = code == 4'hb;
    assign __temp_222 = __reg_state_0 == 6'h37;
    assign __temp_223 = __temp_222 & __temp_221;
    assign __temp_224 = __temp_223 ? 6'h38 : __temp_220;
    assign __temp_225 = code == 4'h3;
    assign __temp_226 = __reg_state_0 == 6'h38;
    assign __temp_227 = __temp_226 & __temp_225;
    assign __temp_228 = __temp_227 ? 6'h39 : __temp_224;
    assign __temp_229 = code == 4'ha;
    assign __temp_230 = __reg_state_0 == 6'h39;
    assign __temp_231 = __temp_230 & __temp_229;
    assign __temp_232 = __temp_231 ? 6'h3a : __temp_228;
    assign __temp_233 = code == 4'hd;
    assign __temp_234 = __reg_state_0 == 6'h3a;
    assign __temp_235 = __temp_234 & __temp_233;
    assign __temp_236 = __temp_235 ? 6'h3b : __temp_232;
    assign __temp_237 = code == 4'he;
    assign __temp_238 = __reg_state_0 == 6'h3b;
    assign __temp_239 = __temp_238 & __temp_237;
    assign __temp_240 = __temp_239 ? 6'h3c : __temp_236;
    assign __temp_241 = code == 4'hd;
    assign __temp_242 = __reg_state_0 == 6'h3c;
    assign __temp_243 = __temp_242 & __temp_241;
    assign __temp_244 = __temp_243 ? 6'h3d : __temp_240;
    assign __temp_245 = code == 4'hb;
    assign __temp_246 = __reg_state_0 == 6'h3d;
    assign __temp_247 = __temp_246 & __temp_245;
    assign __temp_248 = __temp_247 ? 6'h3e : __temp_244;
    assign __temp_249 = code == 4'h4;
    assign __temp_250 = __reg_state_0 == 6'h3e;
    assign __temp_251 = __temp_250 & __temp_249;
    assign __temp_252 = __temp_251 ? 6'h3f : __temp_248;
    assign __reg_state_0_next = __temp_252;

endmodule

